library verilog;
use verilog.vl_types.all;
entity setOnLessThan is
    port(
        inner1          : in     vl_logic_vector(31 downto 0);
        inner2          : in     vl_logic_vector(31 downto 0);
        \out\           : out    vl_logic_vector(31 downto 0)
    );
end setOnLessThan;
