library verilog;
use verilog.vl_types.all;
entity ozer_alican_pr3 is
    port(
        result          : out    vl_logic_vector(31 downto 0)
    );
end ozer_alican_pr3;
