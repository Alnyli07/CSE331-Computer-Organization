library verilog;
use verilog.vl_types.all;
entity test_register is
end test_register;
