library verilog;
use verilog.vl_types.all;
entity test_alu is
end test_alu;
