library verilog;
use verilog.vl_types.all;
entity test_iMem is
end test_iMem;
