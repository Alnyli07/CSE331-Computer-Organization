library verilog;
use verilog.vl_types.all;
entity test_data is
end test_data;
